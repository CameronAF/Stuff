module Mut16_1_test;
reg [15:0] In;
reg [3:0] sel;
wire out;

Mut16_1 M1(out, In, sel);

initial 
begin
	$monitor($time, "out=%b, In=%b, sel=%b\n", out, In, sel);
	#2 In = 16'b0000000000000000; sel = 4'b0000;
	#2 In = 16'b0000000000000001; sel = 4'b0000;
	#2 In = 16'b0000000000000000; sel = 4'b0001;
	#2 In = 16'b0000000000000010; sel = 4'b0001;
	#2 In = 16'b0000000000000000; sel = 4'b0010;
	#2 In = 16'b0000000000000100; sel = 4'b0010;
	#2 In = 16'b0000000000000000; sel = 4'b0011;
	#2 In = 16'b0000000000001000; sel = 4'b0011;
	#2 In = 16'b0000000000000000; sel = 4'b0100;
	#2 In = 16'b0000000000010000; sel = 4'b0100;
	#2 In = 16'b0000000000000000; sel = 4'b0101;
	#2 In = 16'b0000000000100000; sel = 4'b0101;
	#2 In = 16'b0000000000000000; sel = 4'b0110;
	#2 In = 16'b0000000001000000; sel = 4'b0110;
	#2 In = 16'b0000000000000000; sel = 4'b0111;
	#2 In = 16'b0000000010000000; sel = 4'b0111;
	#2 In = 16'b0000000000000000; sel = 4'b1000;
	#2 In = 16'b0000000100000000; sel = 4'b1000;
	#2 In = 16'b0000000000000000; sel = 4'b1001;
	#2 In = 16'b0000001000000000; sel = 4'b1001;
	#2 In = 16'b0000000000000000; sel = 4'b1010;
	#2 In = 16'b0000001000000000; sel = 4'b1010; // this is a repeat In, out will be low
	#2 In = 16'b0000000000000000; sel = 4'b1011;
	#2 In = 16'b0000100000000000; sel = 4'b1011;
	#2 In = 16'b0000000000000000; sel = 4'b1100;
	#2 In = 16'b0001000000000000; sel = 4'b1100;
	#2 In = 16'b0000000000000000; sel = 4'b1101;
	#2 In = 16'b0010000000000000; sel = 4'b1101;
	#2 In = 16'b0000000000000000; sel = 4'b1110;
	#2 In = 16'b0100000000000000; sel = 4'b1110;
	#2 In = 16'b0000000000000000; sel = 4'b1111;
	#2 In = 16'b1000000000000000; sel = 4'b1111;
end
endmodule