/*
 * this module scans the matrix keypad columns with a "walking zero" pattern, 
 * and monitors the keypad rows for a "0" value which indicates that a key has been pressed. 
 * If a "0" is found the column/row value is stored and comapred with the stored value from 
 * the last scan cycle to debounce the keypad. If the column/row value is the same for 2
 * successive scan cycles the keypress is decoded into either a key value (0-9) or 
 * a alaram button (*) or a time button (#) assertion. This block also includes a 
 * key buffer which stores the las 4 keys pressed. New key values are stored in the 
 * buffer when the shift input is pulsed (shift is generated by a FSM block
 * which detects if a new key has been pressed)
*/



module keyscan (clk, reset, shift, rows, columns, key, key_buffer_0, key_buffer_1, key_buffer_2, key_buffer_3, time_button, alarm_button);

input clk, reset, shift;
input [3:0] rows;

output [2:0] columns;
output [3:0] key;
output [3:0] key_buffer_0, key_buffer_1, key_buffer_2, key_buffer_3;
output  time_button, alarm_button;

parameter nokey = 4'b1010;

reg [3:0] new_row, old_row;
reg [2:0] new_column, old_column;

reg [2:0] columns;
reg [3:0] key;
reg [3:0] key_buffer_0, key_buffer_1, key_buffer_2, key_buffer_3;

reg time_button, alarm_button;

always@(posedge clk)
begin
	if(reset)
		columns <=0;
	else
		case (columns)
			3'b111 : columns <= 3'b011;
			3'b011 : columns <= 3'b101;
			3'b101 : columns <= 3'b110;
			3'b110 : columns <= 3'b111;
			default: columns <= 3'b111;
		endcase
end

always@(posedge clk)
begin
	if (reset)
	begin
		new_row <= 0;
		old_row <=0;
		new_column <=0;
		old_column <=0;
		key <= nokey;
		time_button <= 0;
		alarm_button <=0;
	end
	else
	begin
		if (rows[0] == 0 | rows[1] == 0|rows[2] == 0 | rows[3] == 0)
		begin
			new_row <= rows;
			new_column <= columns;
		end
		if(columns == 3'b111)
		begin
			time_button <=0;
			alarm_button <= 0;
			key <= nokey;
			if ((new_row == old_row) & (new_column==old_column))
				case (old_column)
					3'b011:
						case(old_row)
							4'b0111: key <=4'b0001; //1
							4'b1011: key <=4'b0100; //4
							4'b1101: key <=4'b0111; //7
							4'b1110: alarm_button <=1; //* = alarm button
						endcase

					3'b101:
						case(old_row)
							4'b0111: key <=4'b0010; //2
							4'b1011: key <=4'b0101; //5
							4'b1101: key <=4'b1000; //8
							4'b1110: key <=4'b0000; //0
						endcase
					3'b110:
						case(old_row)
							4'b0111: key <=4'b0011; //3
							4'b1011: key <=4'b0110; //6
							4'b1101: key <=4'b1001; //9
							4'b1110: time_button <=1; //# = time button
						endcase
				endcase
				old_row <= new_row;
				old_column <= new_column;
				new_row <= 4'b1111;
				new_column <= 3'b111;
			end
		end
	end
always@(posedge clk)
begin
	if(reset)
	begin
		key_buffer_0 <=0;
		key_buffer_1 <=0;
		key_buffer_2 <=0;
		key_buffer_3 <=0;
	end
	else
		if(shift==1)
		begin
			key_buffer_3 <=key_buffer_2;
			key_buffer_2 <=key_buffer_1;
			key_buffer_1 <=key_buffer_0;
			key_buffer_0 <=key;
		end
end
endmodule