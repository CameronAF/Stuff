module Adder_4bit_test;
reg [3:0] A, B;
wire [4:0] Sum;

Adder_4bit A4bit(Sum, A, B);

initial 
begin
	$monitor($time, "Sum=%b, A=%b, B=%b\n", Sum, A, B);
	#5 A = 4'b0001; B = 4'b0001; //sum = 00010 2
	#5 A = 4'b0101; B = 4'b1110; //sum = 10011 13
	#5 A = 4'b1100; B = 4'b0110; //sum = 10010 12
	#5 A = 4'b1010; B = 4'b0101; //sum = 01111 f
	#5 A = 4'b0101; B = 4'b0010; //sum = 00111 7
	#5 A = 4'b1001; B = 4'b1011; //sum = 10100 14
	#5 A = 4'b0110; B = 4'b0011; //sum = 01001 9
	#5 A = 4'b1111; B = 4'b1111; //sum = 11110 1e
end
endmodule