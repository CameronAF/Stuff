module Adder_4bit(Sum, A, B);
output [4:0] Sum;
input [3:0] A, B;
wire [2:0] C;

HalfAdder HA(Sum[0], C[0], A[0], B[0]);
FullAdder FA1(Sum[1], C[1], A[1], B[1], C[0]);
FullAdder FA2(Sum[2], C[2], A[2], B[2], C[1]);
FullAdder FA3(Sum[3], Sum[4], A[3], B[3], C[2]);
endmodule
